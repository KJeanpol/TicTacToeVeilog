// Verilog testbench code for TIC TAC TOE GAME 

module testbench_Random;

 // Instantiate the Unit Under Test (UUT)
   random ra ();
 // clock

 initial begin
  #100;
  
  #100;
  end
      
endmodule
 