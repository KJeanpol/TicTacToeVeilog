module testbench_Sprite_Controller;
	/*
	logic CLK,
	logic[9:0] x,
	logic[9:0] y,
	logic[7:0] VGA_RED,
	logic[7:0] VGA_GREEN,
	logic[7:0] VGA_BLUE
	
	video_controller UUT (clk, Hsynq, Vsynq, Red, Green, Blue, clk_25Mhz, sync_N, blank_N);
	
	always #5 clk = ~clk;
	*/
	
endmodule
